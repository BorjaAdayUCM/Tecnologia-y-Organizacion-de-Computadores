library IEEE;
use IEEE.STD_LOGIC_1164.all;

package definitions is

	type t_pattern is (no_pattern, first_one, second_one, second_zero, pattern_rec);

end package definitions;